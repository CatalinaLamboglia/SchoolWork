`timescale 1ns/1ps
`include "prj_definition.v"

module mux_tb;
//reg SnA;
//wire CO;//, S;
//wire [31:0] Y;
wire Y;
wire [31:0] Y_32;
wire [31:0] Y_16x1;

reg [31:0] I0_32;
reg [31:0] I1_32;
reg S;
reg I0, I1;

reg [31:0] I0_16x1;
reg [31:0] I1_16x1;
reg [31:0] I2_16x1;
reg [31:0] I3_16x1;
reg [31:0] I4_16x1;
reg [31:0] I5_16x1;
reg [31:0] I6_16x1;
reg [31:0] I7_16x1;
reg [31:0] I8_16x1;
reg [31:0] I9_16x1;
reg [31:0] I10_16x1;
reg [31:0] I11_16x1;
reg [31:0] I12_16x1;
reg [31:0] I13_16x1;
reg [31:0] I14_16x1;
reg [31:0] I15_16x1;

reg [31:0] I16_16x1;
reg [31:0] I17_16x1;
reg [31:0] I18_16x1;
reg [31:0] I19_16x1;
reg [31:0] I20_16x1;
reg [31:0] I21_16x1;
reg [31:0] I22_16x1;
reg [31:0] I23_16x1;
reg [31:0] I24_16x1;
reg [31:0] I25_16x1;
reg [31:0] I26_16x1;
reg [31:0] I27_16x1;
reg [31:0] I28_16x1;
reg [31:0] I29_16x1;
reg [31:0] I30_16x1;
reg [31:0] I31_16x1;

reg [3:0] S_16x1;
reg [4:0] S_32x1;

// module MUX32_2x1(Y, I0, I1, S);
// module MUX1_2x1(Y,I0, I1, S);
MUX1_2x1 mux1(.Y(Y), .I0(I0), .I1(I1), .S(S));
MUX32_2x1 mux2(.Y(Y_32), .I0(I0_32), .I1(I1_32), .S(S));

//MUX32_16x1 mux_16(.Y(Y_16x1), .I0(I0_16x1), .I1(I1_16x1), .I2(I2_16x1), .I3(I3_16x1), .I4(I4_16x1), .I5(I5_16x1),
//               .I6(I6_16x1), .I7(I7_16x1), .I8(I8_16x1), .I9(I9_16x1), .I10(I10_16x1), .I11(I11_16x1),
//               .I12(I12_16x1), .I13(I13_16x1), .I14(I14_16x1), .I15(I15_16x1), .S(S_16x1));

MUX32_32x1 mux_32(.Y(Y_16x1), .I0(I0_16x1), .I1(I1_16x1), .I2(I2_16x1), .I3(I3_16x1), .I4(I4_16x1), .I5(I5_16x1), .I6(I6_16x1), .I7(I7_16x1),
                     .I8(I8_16x1), .I9(I9_16x1), .I10(I10_16x1), .I11(I11_16x1), .I12(I12_16x1), .I13(I13_16x1), .I14(I14_16x1), .I15(I15_16x1),
                     .I16(I16_16x1), .I17(I17_16x1), .I18(I18_16x1), .I19(I19_16x1), .I20(I20_16x1), .I21(I21_16x1), .I22(I22_16x1), .I23(I23_16x1),
                     .I24(I24_16x1), .I25(I25_16x1), .I26(I26_16x1), .I27(I27_16x1), .I28(I28_16x1), .I29(I29_16x1), .I30(I30_16x1), .I31(I31_16x1), .S(S_32x1));


initial 
begin

I0_16x1=0;
I1_16x1=1;
I2_16x1=2;
I3_16x1=3;
I4_16x1=4;
I5_16x1=5;
I6_16x1=6;
I7_16x1=7;
I8_16x1=8;
I9_16x1=9;
I10_16x1=10;
I11_16x1=11;
I12_16x1=12;
I13_16x1=13;
I14_16x1=14;
I15_16x1=15;
I16_16x1=16;
I17_16x1=17;
I18_16x1=18;
I19_16x1=19;
I20_16x1=20;
I21_16x1=21;
I22_16x1=22;
I23_16x1=23;
I24_16x1=24;
I25_16x1=25;
I26_16x1=26;
I27_16x1=27;
I28_16x1=28;
I29_16x1=29;
I30_16x1=30;
I31_16x1=31;

/*#5 ;

I0=1; I1=0; I0_32 = 50; I1_32 = 25; S=0; S_16x1=0;
#5 I0=0; I1=1; I0_32 = 50; I1_32 = 25; S=1; S_16x1=1;
/*#5 S_16x1 = 2 ;
#5 S_16x1 = 3;
#5 S_16x1 = 4 ;
#5 S_16x1 = 5 ;
#5 S_16x1 = 6 ;
#5 S_16x1 = 7 ;
#5 S_16x1 = 8 ;
#5 S_16x1 = 9 ;
#5 S_16x1 = 10 ;
#5 S_16x1 = 11 ;
#5 S_16x1 = 12 ;
#5 S_16x1 = 13 ;
#5 S_16x1 = 14 ;
#5 S_16x1 = 15 ; */
#5 S_32x1 = 0 ;
#5 S_32x1 = 1 ;
#5 S_32x1 = 2 ;
#5 S_32x1 = 3 ;
#5 S_32x1 = 4 ;
#5 S_32x1 = 5 ;
#5 S_32x1 = 6 ;
#5 S_32x1 = 7 ;
#5 S_32x1 = 8 ;
#5 S_32x1 = 9 ;
#5 S_32x1 = 10 ;
#5 S_32x1 = 11 ;
#5 S_32x1 = 12 ;
#5 S_32x1 = 13 ;
#5 S_32x1 = 14 ;
#5 S_32x1 = 15 ;
#5 S_32x1 = 16 ;
#5 S_32x1 = 17 ;
#5 S_32x1 = 18 ;
#5 S_32x1 = 19 ;
#5 S_32x1 = 20 ;
#5 S_32x1 = 21 ;
#5 S_32x1 = 22 ;
#5 S_32x1 = 23 ;
#5 S_32x1 = 24 ;
#5 S_32x1 = 25 ;
#5 S_32x1 = 26 ;
#5 S_32x1 = 27 ;
#5 S_32x1 = 28 ;
#5 S_32x1 = 29 ;
#5 S_32x1 = 30 ;
#5 S_32x1 = 31 ;
end

endmodule